* LMV342 - Rev. A
* Created by Paul Goedeke; April 03, 2019
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2019 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt LMV342 IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID 993F
I_B         22 MID 1P
V_GRp       58 MID 145
V_GRn       59 MID -145
V_ISCp      52 MID 110
V_ISCn      53 MID -110
V_ORn       49 VCLP -2.2
V11         57 48 0
V_ORp       47 VCLP 2.2
V12         56 46 0
V4          41 OUT 0
VCM_MIN     78 VEE_B 0
VCM_MAX     79 VCC_B -600M
I_Q         VCC VEE 70U
XU1         21 22 VOS_DRIFT_0
R69         MID 23 R_NOISELESS 1MEG
GVCCS4      25 MID 24 MID  -167
R63         MID 25 R_NOISELESS 1
R62         MID 24 R_NOISELESS 604K
C21         24 26 26.5F
R61         26 24 R_NOISELESS 100MEG
GVCCS2      26 MID 27 MID  -1
R58         MID 26 R_NOISELESS 1
XCLAWp      VIMON MID 28 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 29 VCCS_LIM_CLAW-_0
R57         MID 27 R_NOISELESS 604K
C16         27 30 26.5F
R56         30 27 R_NOISELESS 100MEG
G_adjust    30 MID ESDp MID  -14.9M
Rsrc        MID 30 R_NOISELESS 1
R55         MID 31 R_NOISELESS 6.5K
C14         31 32 4.9P
R49         32 31 R_NOISELESS 100MEG
GVCCS3      32 MID VCC_B MID  -771M
R48         MID 32 R_NOISELESS 1
R54         MID 33 R_NOISELESS 6.5K
C15         33 34 4.9P
R51         34 33 R_NOISELESS 100MEG
GVCCS1      34 MID VEE_B MID  -771M
R50         MID 34 R_NOISELESS 1
XVCCS_LIM_2 35 MID MID CLAMP VCCS_LIM_2_0
C20         CLAMP MID 13.3N
R94         36 MID R_NOISELESS 1
XZo         37 MID MID 36 VCCS_LIM_ZO_0
R93         37 MID R_NOISELESS 204
C33         37 38 1.59P
R92         37 38 R_NOISELESS 10K
R91         38 MID R_NOISELESS 1
GVCCS11     38 MID 39 MID  -18
C31         40 39 796N
R85         39 MID R_NOISELESS 15.1K
R84         39 40 R_NOISELESS 10K
Rdummy      MID 41 R_NOISELESS 12K
Rx          41 36 R_NOISELESS 120K
R81         40 MID R_NOISELESS 1
GVCCS10     40 MID CL_CLAMP 41  -88.9
Xe_n        ESDp 22 VNSE_0
S5          VEE ESDp VEE ESDp  S_VSWITCH_1
S4          VEE ESDn VEE ESDn  S_VSWITCH_2
S2          ESDn VCC ESDn VCC  S_VSWITCH_3
S3          ESDp VCC ESDp VCC  S_VSWITCH_4
C28         42 MID 1P
R77         43 42 R_NOISELESS 100
C27         44 MID 1P
R76         45 44 R_NOISELESS 100
R75         MID 46 R_NOISELESS 1
GVCCS8      46 MID 47 MID  -1
R74         48 MID R_NOISELESS 1
GVCCS7      48 MID 49 MID  -1
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 22 FEMT_1
GVCCS6      23 MID VSENSE MID  -1U
R68         MID CLAMP R_NOISELESS 1MEG
R44         MID 35 R_NOISELESS 1MEG
XVCCS_LIM_1 50 51 MID 35 VCCS_LIM_1_0
XIQp        VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQn        MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 1P
XCL_AMP     52 53 VIMON MID 54 55 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 56 CLAMP 56  S_VSWITCH_5
SOR_SWn     57 CLAMP 57 CLAMP  S_VSWITCH_6
XGR_AMP     58 59 60 MID 61 62 CLAMP_AMP_HI_0
R39         58 MID R_NOISELESS 1T
R37         59 MID R_NOISELESS 1T
R42         VSENSE 60 R_NOISELESS 1M
C19         60 MID 1F
R38         61 MID R_NOISELESS 1
R36         MID 62 R_NOISELESS 1
R40         61 63 R_NOISELESS 1M
R41         62 64 R_NOISELESS 1M
C17         63 MID 1F
C18         MID 64 1F
XGR_SRC     63 64 CLAMP MID VCCS_LIM_GR_0
R21         54 MID R_NOISELESS 1
R20         MID 55 R_NOISELESS 1
R29         54 65 R_NOISELESS 1M
R30         55 66 R_NOISELESS 1M
C9          65 MID 1F
C8          MID 66 1F
XCL_SRC     65 66 CL_CLAMP MID VCCS_LIM_4_0
R22         52 MID R_NOISELESS 1T
R19         MID 53 R_NOISELESS 1T
R12         28 VCC_B R_NOISELESS 1K
R16         28 67 R_NOISELESS 1M
R13         VEE_B 29 R_NOISELESS 1K
R17         68 29 R_NOISELESS 1M
C6          68 MID 1F
C5          MID 67 1F
G2          VCC_CLP MID 67 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K
G3          VEE_CLP MID 68 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 69 70 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T
R23         VEE_CLP MID R_NOISELESS 1T
R25         69 MID R_NOISELESS 1
R24         MID 70 R_NOISELESS 1
R27         69 71 R_NOISELESS 1M
R28         70 72 R_NOISELESS 1M
C11         71 MID 1F
C10         MID 72 1F
XCLAW_SRC   71 72 CLAW_CLAMP MID VCCS_LIM_3_0
H2          45 MID V11 -1
H3          43 MID V12 1
C12         SW_OL MID 100P
R32         73 SW_OL R_NOISELESS 100
R31         73 MID R_NOISELESS 1
XOL_SENSE   MID 73 44 42 OL_SENSE_0
S1          40 39 SW_OL MID  S_VSWITCH_7
H1          74 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_8
S6          OUT VCC OUT VCC  S_VSWITCH_9
R11         MID 75 R_NOISELESS 1T
R18         75 VOUT_S R_NOISELESS 100
C7          VOUT_S MID 100P
E5          75 MID OUT MID  1
C13         VIMON MID 100P
R33         74 VIMON R_NOISELESS 100
R10         MID 74 R_NOISELESS 1T
R47         76 VCLP R_NOISELESS 100
C24         VCLP MID 100P
E4          76 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K
G8          CLAW_CLAMP MID 23 MID  -1M
R43         MID VSENSE R_NOISELESS 1K
G15         VSENSE MID CLAMP MID  -1M
C4          50 MID 1F
R9          50 77 R_NOISELESS 1M
R7          MID 78 R_NOISELESS 1T
R6          79 MID R_NOISELESS 1T
R8          MID 77 R_NOISELESS 1
XVCM_CLAMP  80 MID 77 MID 79 78 VCCS_EXT_LIM_0
E1          MID 0 81 0  1
R89         VEE_B 0 R_NOISELESS 1
R5          82 VEE_B R_NOISELESS 1M
C3          82 0 1F
R60         81 82 R_NOISELESS 1MEG
C1          81 0 1
R3          81 0 R_NOISELESS 1T
R59         83 81 R_NOISELESS 1MEG
C2          83 0 1F
R4          VCC_B 83 R_NOISELESS 1M
R88         VCC_B 0 R_NOISELESS 1
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       84 80 R_NOISELESS 1K
G_PSR       80 84 31 33  -1M
R2          51 ESDn R_NOISELESS 1M
R1          84 85 R_NOISELESS 1M
R_CMR       21 85 R_NOISELESS 1K
G_CMR       85 21 25 MID  -1M
C_CMn       ESDn MID 5P
C_CMp       MID ESDp 5P
R53         ESDn MID R_NOISELESS 1T
R52         MID ESDp R_NOISELESS 1T
R35         IN- ESDn R_NOISELESS 10M
R34         IN+ ESDp R_NOISELESS 10M

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_8 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_9 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)

.ENDS LMV342
*
.SUBCKT VOS_DRIFT_0  VOS+ VOS-
.PARAM DC = 25U
.PARAM POL = -1
.PARAM DRIFT = 1.9E-6
E1 VOS+ VOS- VALUE={DC+POL*DRIFT*(TEMP-27)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0.05351, 1.01E-06)
+(1.5108, 2.39E-05)
+(11.723, 1.85E-04)
+(52.59, 8.82E-04)
+(80.92, 1.55E-03)
+(105.11, 2.60E-03)
+(106.38, 2.75E-03)
+(124.67, 4.90E-03)
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0.0382, 1.11E-06)
+(10.233, 2.53E-04)
+(60.300, 1.69E-03)
+(85.760, 2.749E-03)
.ENDS
*


.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 2.54E-3
.PARAM IPOS = 1.52E-2
.PARAM INEG = -1.52E-2
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 5
.PARAM IPOS = 28K
.PARAM INEG = -28K
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=190
.PARAM NVR=24
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=24
.PARAM NVRF=24
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT FEMT_1  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=1
.PARAM NVRF=1
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 4
.PARAM INEG = -4
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.9
.PARAM INEG = -0.9
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.35
.PARAM INEG = -0.35
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*


